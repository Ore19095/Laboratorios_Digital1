module testbench();
    reg D1,D0;
    reg S0;
    wire out;

endmodule